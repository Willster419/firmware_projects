/////////////////////////////////////////////////////////////////////
// pipeline_tb.sv
// simple device testbench
// Willster419
// 2020/07/31
// A simple testbench for simulating the pipeline module
/////////////////////////////////////////////////////////////////////
