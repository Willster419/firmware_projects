---------------------------------------------------------------------
-- hello_world.vhd
-- top design module
-- Willster419
-- 2020-07-31
-- 
---------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity hello_world is
  generic (

  );
  port (
    
  );
end entity hello_world;

architecture rtl of hello_world is
  
begin
  
  
  
end architecture hello_world;
