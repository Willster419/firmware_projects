---------------------------------------------------------------------
-- hello_world.vhd
-- top design module
-- Willster419
-- 2020-07-31
-- A pipeline module for adding delay to a sample design
---------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pipeline is
  generic (

  );
  port (
    
  );
end entity pipeline;

architecture rtl of pipeline is
  
begin
  
  
  
end architecture rtl;
